library verilog;
use verilog.vl_types.all;
entity moving_average_filter_vlg_vec_tst is
end moving_average_filter_vlg_vec_tst;
